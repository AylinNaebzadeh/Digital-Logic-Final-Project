--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   10:57:45 01/13/2022
-- Design Name:   
-- Module Name:   D:/Logical-Circute/Final-Project-VHDL/secondTry/Counter_tb.vhd
-- Project Name:  secondTry
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: Counter
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY Counter_tb IS
END Counter_tb;
 
ARCHITECTURE behavior OF Counter_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT Counter
    PORT(
         CLK : IN  std_logic;
         RST : IN  std_logic;
         COUNT : INOUT  std_logic_vector(4 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal CLK : std_logic := '1';
   signal RST : std_logic := '1';

	--BiDirs
   signal COUNT : std_logic_vector(4 downto 0);

   -- Clock period definitions(it has been commented by me)
   --constant CLK_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: Counter PORT MAP (
          CLK => CLK,
          RST => RST,
          COUNT => COUNT
        );

   -- Clock process definitions
   CLK_process :process
   begin
		RST <= '0';
		CLK <= '0';
		wait for 20 ns;
		CLK <= '1';
   end process;
 

   -- Stimulus process
   --stim_proc: process
   --begin		
      -- hold reset state for 100 ns.
      --wait for 100 ns;	

      --wait for CLK_period*10;

      -- insert stimulus here 

      --wait;
   --end process;

END;
